// Test file for Verilog parser

module test_module(input a, input b, output c, output d, wire e, reg f);
endmodule
