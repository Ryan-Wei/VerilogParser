// comment0
// comment1


module test_module(input a, input b, output c, output d, wire e, reg f); // uycucyc
    reg x;
    input [4:0] y;
    always @ (x)
    begin
        if(x)
            yyy;
        else
            zzz;
    end
    always @ (2)
    begin
        yyyyy;
        begin
            1+1;
            zzzzz;
            if (xixi)
            begin
                haha;
                hehe;
            end
        end
    end


endmodule

//module ALU(w,t,c,s,reg [0:3] y); // uycucyc
//endmodule